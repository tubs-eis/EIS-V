library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library eisv;
use eisv.eisv_types_pkg.all;

entity eisv_ctrl is
    port (
        instruction_i : in decoded_instruction_t;
        ctrl_o : out control_word_t
    );
end entity;

architecture gen of eisv_ctrl is

    type ctrl_table_t is array (0 to 2047) of control_word_t;

    constant CTRL_TABLE : ctrl_table_t := (
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ZERO, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '1', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', SHIFTER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', SHIFTER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, NOT_ZERO, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', OP_A, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', WORD, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', CONDITION, '1', EXECUTION_UNIT, REG, IMM, '1', '0', '^', LEFT, MUL, DIV, LESS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', WORD, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', CONDITION, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, LESS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', CONDITION, '1', EXECUTION_UNIT, REG, IMM, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', CONDITION, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', CLEAR, LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '1', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, LESS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', SHIFTER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', RIGHT_LOGICAL, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', SHIFTER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', RIGHT_LOGICAL, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_LESS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', OP_A, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '&', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '&', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, CARRY, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', CLEAR, LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ZERO, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '1', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', SHIFTER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', SHIFTER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, NOT_ZERO, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', OP_A, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', WORD, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', CONDITION, '1', EXECUTION_UNIT, REG, IMM, '1', '0', '^', LEFT, MUL, DIV, LESS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', WORD, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', CONDITION, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, LESS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', CONDITION, '1', EXECUTION_UNIT, REG, IMM, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', CONDITION, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', CLEAR, LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '1', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, LESS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', HALF, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', SHIFTER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', RIGHT_ARITHMETIC, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', SHIFTER, '1', EXECUTION_UNIT, REG, REG, '0', '0', '^', RIGHT_ARITHMETIC, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_LESS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', OP_A, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, NOT_CARRY, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', '|', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '1', '0', '1', '0', ADDER, '0', LOAD_STORE_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', LOGIC, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '&', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, PC, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '1', '1', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, REG, REG, '0', '0', '&', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, REG, REG, '1', '0', '^', LEFT, MUL, DIV, CARRY, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '1', '0', ADDER, '1', PC_PLUS_4, REG, IMM, '0', '1', '^', LEFT, MUL, DIV, ALWAYS, '1', EU_RESULT, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '1', '1', '0', '0', '0', ADDER, '1', PC_PLUS_4, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '1', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', LOGIC, '1', EXECUTION_UNIT, RS1, IMM, '0', '0', CLEAR, LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '1', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' ),
        ( '0', '0', '0', '1', '1', ADDER, '1', EXECUTION_UNIT, ZERO, IMM, '0', '0', '^', LEFT, MUL, DIV, ALWAYS, '0', PC_OFFSET, '0', '0', BYTE, '0', '0', '0', '0', '0', '0', UNIMPLEMENTED, MEPC, '0', '0', '0' )
    );
begin

    decode: process (all) is
        variable control_bits : unsigned(10 downto 0);
    begin
        control_bits := instruction_i.funct7(5) & instruction_i.funct3(2) & instruction_i.funct3(1) & instruction_i.funct3(0) & instruction_i.opcode(6) & instruction_i.opcode(5) & instruction_i.opcode(4) & instruction_i.opcode(3) & instruction_i.opcode(2) & instruction_i.opcode(1) & instruction_i.opcode(0);
        ctrl_o <= CTRL_TABLE(to_integer(unsigned(control_bits)));
    end process;

end architecture;
